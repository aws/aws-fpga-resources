version https://git-lfs.github.com/spec/v1
oid sha256:7d5a195679e89f11e020d2ee65f4348cf407cb50aa4fc1e806b39c0700849cc8
size 6064
