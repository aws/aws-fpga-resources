version https://git-lfs.github.com/spec/v1
oid sha256:b5b15e256ddc2d95b22ffbfd63d1eee418ea6fc0edd50577f65db14d3bd20fd3
size 17474
