version https://git-lfs.github.com/spec/v1
oid sha256:a91b5275dc0ad30bea4cb44779468700c3ac010471b80c16ee42809223824d10
size 5820
