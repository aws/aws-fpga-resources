version https://git-lfs.github.com/spec/v1
oid sha256:76706521177b92af73b5cd639c7c2e0a14e1325deca5258a270eeb571054c8e9
size 6073
