version https://git-lfs.github.com/spec/v1
oid sha256:d24c96458d399a50caa06068d2d74827dd5bc8b540c33761de7f7c9409537be9
size 6065
