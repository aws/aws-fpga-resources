version https://git-lfs.github.com/spec/v1
oid sha256:7d45a70f745c5f3da7b71d23c66158d5cc3cf6abbd74e8f75e46547858e9267b
size 6065
