version https://git-lfs.github.com/spec/v1
oid sha256:7f31713aa566b74eff78bfc2a52f0ecc26682745fd5176a8ac47df167e0401fc
size 6944
