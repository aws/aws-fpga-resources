version https://git-lfs.github.com/spec/v1
oid sha256:74bce4abbcdfcf693e51755e6ab710b0b63a7a7b96611d2e5d57b5d4f9122171
size 6323
