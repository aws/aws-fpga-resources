version https://git-lfs.github.com/spec/v1
oid sha256:66a8bdfc8275be11f472b910ba809cf8abe0b5a7337f5122c09805f8ec8651fe
size 6932
