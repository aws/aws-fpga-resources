version https://git-lfs.github.com/spec/v1
oid sha256:12862bf8fc4e93c1799652cc0dc22745603ac11eb41aaf2f2de5580a8b061613
size 286032
