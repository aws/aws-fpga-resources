version https://git-lfs.github.com/spec/v1
oid sha256:b0152d8f81a01b384a4640a878b33761921f0e86d3a62fdcfbce1d24db9db324
size 6322
