version https://git-lfs.github.com/spec/v1
oid sha256:8c3120c1a0722bc5a14970e9a7f953142c991f27636800823cf5e1af0f99dc31
size 13220
