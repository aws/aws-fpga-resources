version https://git-lfs.github.com/spec/v1
oid sha256:0cbf88c90ddf6bc0cff5b10d5198ea984f008a1af4fd25d552599a54c0898e7e
size 248055
