version https://git-lfs.github.com/spec/v1
oid sha256:a1099b55da62c2bab9726141526a40eed24e614a7459a235fcf7e510c7a2a4d3
size 334315
