version https://git-lfs.github.com/spec/v1
oid sha256:4417b94ff2f288698d0b808b8c9fff3bba5d5bf3eacd54b046ebce8026324fc0
size 7669
