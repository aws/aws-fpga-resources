version https://git-lfs.github.com/spec/v1
oid sha256:8c06592df94920cb8305c0b39ef89e4cb49c4d4e9f1c93aece0a3f63888b7056
size 416774
