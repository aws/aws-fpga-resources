version https://git-lfs.github.com/spec/v1
oid sha256:611fa548ddd4a750692d27429cb850a8ece19b0b3ad91712aad535721ffcf235
size 6075
