version https://git-lfs.github.com/spec/v1
oid sha256:00da2c392aa76b9ef3a63b7e752e9b46ad0165bac757ed91341b6cd4e32b5ac2
size 13229
