version https://git-lfs.github.com/spec/v1
oid sha256:cfc8714fa2c9b81dce16ddb6c2aa23611cd150da47e2ca1099af9b027ce07c35
size 18419
