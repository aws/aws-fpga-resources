version https://git-lfs.github.com/spec/v1
oid sha256:860a6153a890bf9018156595e322b40f4df768624c0a2126357f5a53a5cb9c4d
size 6066
