version https://git-lfs.github.com/spec/v1
oid sha256:e619b3e05c0730b43465c5c750be5bee489d1ff418027bc33e2ed17f5ec7d5ec
size 7419
