version https://git-lfs.github.com/spec/v1
oid sha256:c61d4473d93631ab617450fcff57d468895238e8626421c416980718461df823
size 6943
