version https://git-lfs.github.com/spec/v1
oid sha256:a6fc9efd90b4c30ca9731c16f73670975f44c06f707b90eb898679dc9a99bd69
size 17009
