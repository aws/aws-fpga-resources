version https://git-lfs.github.com/spec/v1
oid sha256:7b75a051bc74ed753154bf7c875203e0eaa2d8cb52466d7b1a872bda42a7221c
size 6962
