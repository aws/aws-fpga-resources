version https://git-lfs.github.com/spec/v1
oid sha256:fa41b6cb23b7c373657b3b0c2cef1ba0d2d303f02964ccb50825131585bb197d
size 7413
