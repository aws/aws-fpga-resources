version https://git-lfs.github.com/spec/v1
oid sha256:7d74e166a0cc8a3d4c62d5cf73feb8a376dc3289f50d97b1f1b87009401c1801
size 7669
