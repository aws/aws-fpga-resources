version https://git-lfs.github.com/spec/v1
oid sha256:ca5258befb31609b14197ec9435dd495b5abcb4d787bbb7ff5b2daa51563d1e1
size 6786
