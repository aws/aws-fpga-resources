version https://git-lfs.github.com/spec/v1
oid sha256:98e1a439d52859140723e5f6e1c9ee590d48a7900a67cf1b1ccdb8701c6153d1
size 15998
