version https://git-lfs.github.com/spec/v1
oid sha256:e4663829b76b8642985fb91686b7812c4b19f913bbbeb1acc47615eb92d9bbbf
size 6954
