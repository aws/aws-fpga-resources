version https://git-lfs.github.com/spec/v1
oid sha256:b87b5e8ebb73c4d4ce32e233bd104b3213017c034a6bd89ea457a5c37652b38f
size 17214
