version https://git-lfs.github.com/spec/v1
oid sha256:2cf9cd58f6f48514740cf9eb2426bad544e9d7c4775ef122a73ef2e985215a08
size 7389
