version https://git-lfs.github.com/spec/v1
oid sha256:2441edcfcf3717a754e1239dc04d963a9bf2cd6adb1d092a740b4b239c93a800
size 26922
