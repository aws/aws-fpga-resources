version https://git-lfs.github.com/spec/v1
oid sha256:c9989d5ddccac5bfcfefcc86f09e1351478ac6b492f77e95633c2e342e15ed43
size 16004
