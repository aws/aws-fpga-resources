version https://git-lfs.github.com/spec/v1
oid sha256:8dce457abf3f8ddf06ea1477ad227f0602f9fac3bbfd38e7483c49178ccd9e05
size 17514
