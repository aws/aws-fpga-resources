version https://git-lfs.github.com/spec/v1
oid sha256:2feef6be118f58b24c915caf86659a52856ed296a8b02f642661e05678f2e744
size 6064
