version https://git-lfs.github.com/spec/v1
oid sha256:c891d07012de0702aad878621b3bfadae1caa30fc99ec464bc01ac0fbc303e03
size 31032
