version https://git-lfs.github.com/spec/v1
oid sha256:92411fc22ee7a42fbf2659aa518ab6827dcb121371559389d342089887ddbae5
size 18069
