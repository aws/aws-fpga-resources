version https://git-lfs.github.com/spec/v1
oid sha256:283b639b26900cc0c6c92df0477625b93137574a0f9a96f81f251b01aa3c391a
size 16970
