version https://git-lfs.github.com/spec/v1
oid sha256:3df952b4fb8d65b54699f395fa6b32fa3c185d2c9c89a54e524f01bf114d3082
size 6067
