version https://git-lfs.github.com/spec/v1
oid sha256:6410f0463e98c7dff1a7716f1ec45ecdf80b4acf41cc034dac6045bb6a0fc0dc
size 17277
