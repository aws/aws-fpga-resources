version https://git-lfs.github.com/spec/v1
oid sha256:2774a06132b3237cbefd9217bfee4fc92e5007c1c5bc3664d3f6edf1fa8919fb
size 6073
