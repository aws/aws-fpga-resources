version https://git-lfs.github.com/spec/v1
oid sha256:958dfa1c811cfafa92edf3c72f69ddbc389e643558f9df0c76aadc6d74af447c
size 13979
