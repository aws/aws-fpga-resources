version https://git-lfs.github.com/spec/v1
oid sha256:d84dd8339d73ca3718a3167c5d919d0374e6ced17b0d41873a7105cb05b30ad9
size 18344
