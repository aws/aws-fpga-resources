version https://git-lfs.github.com/spec/v1
oid sha256:d5d5ed4d02e9ef160cc3adb49597e3019ed5c176fbd786473c5c3cb7faa052a4
size 16004
