version https://git-lfs.github.com/spec/v1
oid sha256:28c8fc04f86d320a7487be2fa957852f1acb35dcf7e8ba9f5779e01534687053
size 7678
