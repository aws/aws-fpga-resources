version https://git-lfs.github.com/spec/v1
oid sha256:5e0454beb355f5c2ecd2451ef98f73fb8e183951042f68a2244aa724d61b2fe1
size 6067
