version https://git-lfs.github.com/spec/v1
oid sha256:bcc679cc6f43ab4483f564a2efc9bf7a2991493b9a4620fe27a2143dcf30f0aa
size 13229
