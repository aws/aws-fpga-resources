version https://git-lfs.github.com/spec/v1
oid sha256:45b0c501d78e433e9b875dedd4b779b8b61175b78de2aae4ce9adf43aea70b02
size 7678
