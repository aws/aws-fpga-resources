version https://git-lfs.github.com/spec/v1
oid sha256:e4598c709a8532c9f3276cad4ab0e377f9877dffcf633601ba0ce24fde4b99d4
size 6960
