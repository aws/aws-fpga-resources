version https://git-lfs.github.com/spec/v1
oid sha256:d2eef8e6d72e58e23709b391b39c8f86a8942c8fb2d9e077201d78fd14acc9f6
size 5797
