version https://git-lfs.github.com/spec/v1
oid sha256:64ff2ed60e1ecc9e62fa4fe6245d29457a55c694f86ee6421582dfc3f5b5afda
size 13970
