version https://git-lfs.github.com/spec/v1
oid sha256:e0928b541da4e3369311c7a99afd9f6bdd6c5b4a05353eabac80fe77dc670bcc
size 6072
