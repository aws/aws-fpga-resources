version https://git-lfs.github.com/spec/v1
oid sha256:67d8dd425bf8a226257bf427607e8c78854f6725e5750988aa4ded1da5a304f9
size 6943
