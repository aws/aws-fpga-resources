version https://git-lfs.github.com/spec/v1
oid sha256:bc1b8629468527aff17bd4169f1d4ec9ae862cee70eb49bd4a8c66533b61bace
size 6779
