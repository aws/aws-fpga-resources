version https://git-lfs.github.com/spec/v1
oid sha256:ddefda593132528604d17f576de9fc4d12c3a74d209d79d0d7d91e837e25061a
size 6072
