version https://git-lfs.github.com/spec/v1
oid sha256:068774d0009a328fdd2e9d72e4a5379282e3f9eef8a4a93625af4e9a8e21ec68
size 6074
