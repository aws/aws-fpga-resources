version https://git-lfs.github.com/spec/v1
oid sha256:b69de831e7624dc337b9cc4e4c60280802d9f300ed9c88ae7c51204f8728be28
size 17263
