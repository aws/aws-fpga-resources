version https://git-lfs.github.com/spec/v1
oid sha256:c003b06359902b377b8f8d45d22ed4b789e55b190621128dd4a4e84cfab158cc
size 6323
