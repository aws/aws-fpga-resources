version https://git-lfs.github.com/spec/v1
oid sha256:f46ced075743e958f9ff20b305d935b02b3b0e494d98f37ad911a5f340e6d589
size 6075
