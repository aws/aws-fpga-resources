version https://git-lfs.github.com/spec/v1
oid sha256:d2264499a4743d2745ed489e504a59d7bec1c5b094881e9c4fdf3fd74aa3ee4e
size 13970
