version https://git-lfs.github.com/spec/v1
oid sha256:bcd4e57252ab5ec472dd1a6671e7de58a096504620943e46c609631f82a614a2
size 8225
