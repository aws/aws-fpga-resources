version https://git-lfs.github.com/spec/v1
oid sha256:2b6916723b071ba8303df9ccfc6e7fb176bcd4e3e5f6dcd578ba65be75e56ac9
size 6057
