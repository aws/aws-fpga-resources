version https://git-lfs.github.com/spec/v1
oid sha256:b1f4154be5fd076443647b90bd7ac8956107edc0881909a5023dc9b11023b1a8
size 6074
