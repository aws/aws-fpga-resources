version https://git-lfs.github.com/spec/v1
oid sha256:7a6e29617234da55dc909d3dadefa6a060ac330d17c6a5edaba557e938be5771
size 13229
