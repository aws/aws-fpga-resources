version https://git-lfs.github.com/spec/v1
oid sha256:8f954e87ac9247cef92bd478c262eeb08a5eb06b1126dbbc3727aee0153820c8
size 13220
