version https://git-lfs.github.com/spec/v1
oid sha256:8cd49e7de36287557d87a4f005f905c5dbf692a30c1978afe34088317e369ca1
size 17514
