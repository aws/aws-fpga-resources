version https://git-lfs.github.com/spec/v1
oid sha256:0507d9ccf0d8a3d6f0e238d6607e52d8945908d13bffb5f150f2d3b704546381
size 17009
