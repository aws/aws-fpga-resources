version https://git-lfs.github.com/spec/v1
oid sha256:a30eaa11e63139651682ded698a5d9f64ffd9121e2e95302583e6bb310cc8411
size 8214
