version https://git-lfs.github.com/spec/v1
oid sha256:b76e41370268e8f44ab32e2d27d4910268f5be51ccf5bfe2f94f711f2cce93dd
size 18381
