version https://git-lfs.github.com/spec/v1
oid sha256:85c104eb322683a0602bbe3b355b171f874c6f66ec81ffab617c1aaeead80604
size 18419
