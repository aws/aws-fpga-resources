version https://git-lfs.github.com/spec/v1
oid sha256:3c152011ab6a8be7790a128c3828ec4ad4624d9113b087bd778732dc09d74ecb
size 6962
