version https://git-lfs.github.com/spec/v1
oid sha256:1c887e460726a2fcbdc0bb65a49ff38b0b8912c9155a7719f41043ba4a386972
size 16995
