version https://git-lfs.github.com/spec/v1
oid sha256:c047b2a75486a7bd3f4a68397d12373905f69b7cbc77da6214f3fc00790ea5bf
size 6072
