version https://git-lfs.github.com/spec/v1
oid sha256:5e38e2ca19c4bd58ba28fcef336a48fcb91b3edf4d999f81fe1811bbddfb31db
size 17514
