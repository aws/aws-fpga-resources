version https://git-lfs.github.com/spec/v1
oid sha256:b303a499c58b665c369556f33830789009dc319c0348d0f2db0be77bf241516a
size 6066
