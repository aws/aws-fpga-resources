version https://git-lfs.github.com/spec/v1
oid sha256:c549b1bccd470935e9d20a7e161f9f433679427ab22cabb4a5b9a745a0c0149f
size 6072
