version https://git-lfs.github.com/spec/v1
oid sha256:99fe99b6b5911a2a1ebbc65a9a0844f788bb3849d38b431fa94b58163010dc5d
size 18381
