version https://git-lfs.github.com/spec/v1
oid sha256:f058df8f68a1e36638b2aa73707e46a9cdb530595998695045be1a50c10737b9
size 6950
