version https://git-lfs.github.com/spec/v1
oid sha256:78ba2a06833d3c35bb8fa35cdcc9e4c6a4a0cef5d346a4010b701edb4d962366
size 7413
