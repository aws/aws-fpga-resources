version https://git-lfs.github.com/spec/v1
oid sha256:70e0574a473bebe221544796fff4c8aa56d896342a2967d9c5197429cd36d38f
size 6959
