version https://git-lfs.github.com/spec/v1
oid sha256:736cf64d3cc850a3f4c66d610459f4dd1f9c5f65fe4916ceee88f72820127315
size 13979
