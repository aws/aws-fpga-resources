version https://git-lfs.github.com/spec/v1
oid sha256:752fb995904d528ca7abb51cefa06102ea5e19050f847cd92b8f88dc65c8819d
size 6954
