version https://git-lfs.github.com/spec/v1
oid sha256:8830ba3288d06fbc8014cf98f658fb3ceee7d2083ff1680ddb5efdd43c5cd2e6
size 8170
