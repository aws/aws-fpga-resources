version https://git-lfs.github.com/spec/v1
oid sha256:af0b875fbb47221d730287ac358389a7aa4004f3d958d428853bda86d152bfac
size 3246093
