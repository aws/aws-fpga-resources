version https://git-lfs.github.com/spec/v1
oid sha256:48e38d4a2ef24164e0270ace048e512b32a9c43b07cda70a582468083ae731a0
size 18283
