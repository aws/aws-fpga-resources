version https://git-lfs.github.com/spec/v1
oid sha256:8055b7af5724f92f1af0b3e9dbdd086152019c55f5eac396e440372acf4fed75
size 6944
