version https://git-lfs.github.com/spec/v1
oid sha256:dd735739b4f3ccc298635afc04739b5cf4130598e4d0043ce35ead9bef5083b6
size 5820
