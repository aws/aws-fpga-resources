version https://git-lfs.github.com/spec/v1
oid sha256:0fed48d26d5603052a6fa3163a1a43c99d9f874a2f258942a246492832286dcb
size 6962
