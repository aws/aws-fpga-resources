version https://git-lfs.github.com/spec/v1
oid sha256:e867f4485f32531bf72a5821aa7e7f34dff829be31b847154bd1f35f8bbf7a0d
size 18344
