version https://git-lfs.github.com/spec/v1
oid sha256:8440cd52e50cc4777d7d72426bd93b2fc3a97cba88f3332c770e5e0060fbfa55
size 6967
