version https://git-lfs.github.com/spec/v1
oid sha256:d7f1b5b6af83cbfa0bdb436d6608a6b39313ef21b05c2d4467be29d3c7ed0244
size 13220
