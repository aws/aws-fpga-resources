version https://git-lfs.github.com/spec/v1
oid sha256:0396b0276be858d6f1ef6618446bfbf74d82da814763cf9a6b07604cdbe8c60b
size 6960
