version https://git-lfs.github.com/spec/v1
oid sha256:33f0b555cc868c82072abc8a4eaf0f60bdf1e7ee49bf6f6f265a75451c31ecb7
size 6786
