version https://git-lfs.github.com/spec/v1
oid sha256:0b575a23f8c134a099dd3b0a0d4db090f9b5ceb1db13033bb42ee4c48c29c1dc
size 17263
