version https://git-lfs.github.com/spec/v1
oid sha256:f1cf69807fc445613f84dd328fa7b267853739041f81615bcb8955f6cc20ee0e
size 6295
