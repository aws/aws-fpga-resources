version https://git-lfs.github.com/spec/v1
oid sha256:979a4f196ba3e7009955b99a53e51b67a9a3921e191f4b9250fa4363363a9800
size 6959
