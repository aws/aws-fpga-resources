version https://git-lfs.github.com/spec/v1
oid sha256:2ec34bd516df12fc729bcd4b31b00ad841556f8e32b2a24ff7863862dcb80d51
size 6959
