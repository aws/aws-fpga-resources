version https://git-lfs.github.com/spec/v1
oid sha256:94840c0410ad69ffde6ba1a2d3c345e8aec7ea8a8db60212ec0ca1acbd2c15b2
size 67896
