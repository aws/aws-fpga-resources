version https://git-lfs.github.com/spec/v1
oid sha256:eb012651a1e27813a473beb7fdd3cc30945ecba799d481ae33364809b5c7dd7e
size 6959
