version https://git-lfs.github.com/spec/v1
oid sha256:24231c8a3e179aeed960afac99b1f538a9dc31cf07a9c8ae9cd15b534d5d0731
size 111192
