version https://git-lfs.github.com/spec/v1
oid sha256:0959f72c2f5681092bac387b1dd48547fdd8ba6381db866ac4bb8db160e85afa
size 6950
