version https://git-lfs.github.com/spec/v1
oid sha256:40dbe316383d2ed2571045ca7b6d85c31d9dba485c52ef4d6e701674fb93483e
size 6073
