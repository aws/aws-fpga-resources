version https://git-lfs.github.com/spec/v1
oid sha256:b1faceac085b3025483512b698ac2263bad79a56c1b19e68bd85a273359df991
size 26942
