version https://git-lfs.github.com/spec/v1
oid sha256:0f62b9a9d4b2843f9488e8aa865d86b4da45000495b44c185756a70cefdeacc2
size 13970
