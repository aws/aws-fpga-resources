version https://git-lfs.github.com/spec/v1
oid sha256:33527029a081f095fa1307e50fe9e77dc133fe532804d70d45cd73080bd2a80e
size 6962
