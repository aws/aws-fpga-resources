version https://git-lfs.github.com/spec/v1
oid sha256:c59dec456605375a7bfd7e60036830f5c5b87d37f797aa76ebaa32b69d4ce171
size 6322
