version https://git-lfs.github.com/spec/v1
oid sha256:6afea3f9a3dade0732bde2054afd01be7b7a7afeec26c905d4fa9278933e7d5a
size 6967
