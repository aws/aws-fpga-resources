version https://git-lfs.github.com/spec/v1
oid sha256:c262b26cd2412b9a1d1ef8a79e8d1d64d4dd093d7544e1de2475f6f87a4c251f
size 86188
