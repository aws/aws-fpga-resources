version https://git-lfs.github.com/spec/v1
oid sha256:fa67fb29b8d4d2117b41d124ce731d7adb55f59d21217ea8a98e5eb299ca6b04
size 8214
