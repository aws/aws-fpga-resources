version https://git-lfs.github.com/spec/v1
oid sha256:b4b6dea1d122a106bf04a1857f0b52afb2ee60a595343198b4ef6facae0568fc
size 5823
