version https://git-lfs.github.com/spec/v1
oid sha256:3d46556ce65cfb61c7e5218db522e5ba021879cce8f178b6dc7751b400742052
size 5823
