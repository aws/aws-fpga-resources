version https://git-lfs.github.com/spec/v1
oid sha256:348df2cc40299c0095fc7b82729058d853701bb3b924c3b5d52bda84bf555fc0
size 6073
