version https://git-lfs.github.com/spec/v1
oid sha256:5efccab062244d7cfacc6beb187e488ac2a66c995a3ff02886408dc707fea5b7
size 18344
