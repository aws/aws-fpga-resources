version https://git-lfs.github.com/spec/v1
oid sha256:1ba275648f8d1f0b571b9bd4ab54755b0f447877f70f1682d09d542222c6768b
size 13979
