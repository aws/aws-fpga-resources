version https://git-lfs.github.com/spec/v1
oid sha256:6ce7f252c96550cf73a0c4795b3426463819f87f45b232774b4083a50cec20c7
size 17277
