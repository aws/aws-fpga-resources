version https://git-lfs.github.com/spec/v1
oid sha256:4e58a3da1bd397fe34a090432d9092b7c3f04891ce79374f776c2c3c68e88573
size 6779
